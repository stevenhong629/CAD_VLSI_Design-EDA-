`timescale 1ns/1ps
module c880 (gat1, gat8, gat13, gat17, gat26, gat29, gat36, gat42, gat51, gat55, gat59, gat68, gat72, gat73, gat74, gat75, gat80, gat85, gat86, gat87, gat88, gat89, gat90, gat91, gat96, gat101, gat106, gat111, gat116, gat121, gat126, gat130, gat135, gat138, gat143, gat146, gat149, gat152, gat153, gat156, gat159, gat165, gat171, gat177, gat183, gat189, gat195, gat201, gat207, gat210, gat219, gat228, gat237, gat246, gat255, gat259, gat260, gat261, gat267, gat268, gat_out388, gat_out389, gat_out390, gat_out391, gat_out418, gat_out419, gat_out420, gat_out421, gat_out422, gat_out423, gat_out446, gat_out447, gat_out448, gat_out449, gat_out450, gat_out767, gat_out768, gat_out850, gat_out863, gat_out864, gat_out865, gat_out866, gat_out874, gat_out878, gat_out879, gat_out880);
input gat1, gat8, gat13, gat17, gat26, gat29, gat36, gat42, gat51, gat55, gat59, gat68, gat72, gat73, gat74, gat75, gat80, gat85, gat86, gat87, gat88, gat89, gat90, gat91, gat96, gat101, gat106, gat111, gat116, gat121, gat126, gat130, gat135, gat138, gat143, gat146, gat149, gat152, gat153, gat156, gat159, gat165, gat171, gat177, gat183, gat189, gat195, gat201, gat207, gat210, gat219, gat228, gat237, gat246, gat255, gat259, gat260, gat261, gat267, gat268;
output gat_out388, gat_out389, gat_out390, gat_out391, gat_out418, gat_out419, gat_out420, gat_out421, gat_out422, gat_out423, gat_out446, gat_out447, gat_out448, gat_out449, gat_out450, gat_out767, gat_out768, gat_out850, gat_out863, gat_out864, gat_out865, gat_out866, gat_out874, gat_out878, gat_out879, gat_out880;
wire gat_out269, gat_out270, gat_out273, gat_out276, gat_out279, gat_out280, gat_out284, gat_out285, gat_out286, gat_out287, gat_out290, gat_out291, gat_out292, gat_out293, gat_out294, gat_out295, gat_out296, gat_out297, gat_out298, gat_out301, gat_out302, gat_out303, gat_out304, gat_out305, gat_out306, gat_out307, gat_out308, gat_out309, gat_out310, gat_out316, gat_out317, gat_out318, gat_out319, gat_out322, gat_out323, gat_out324, gat_out325, gat_out326, gat_out327, gat_out328, gat_out329, gat_out330, gat_out331, gat_out332, gat_out333, gat_out334, gat_out335, gat_out336, gat_out337, gat_out338, gat_out339, gat_out340, gat_out341, gat_out342, gat_out343, gat_out344, gat_out345, gat_out346, gat_out347, gat_out348, gat_out349, gat_out350, gat_out351, gat_out352, gat_out353, gat_out354, gat_out355, gat_out356, gat_out357, gat_out360, gat_out363, gat_out366, gat_out369, gat_out375, gat_out376, gat_out379, gat_out382, gat_out385, gat_out392, gat_out393, gat_out399, gat_out400, gat_out401, gat_out402, gat_out403, gat_out404, gat_out405, gat_out406, gat_out407, gat_out408, gat_out409, gat_out410, gat_out411, gat_out412, gat_out413, gat_out414, gat_out415, gat_out416, gat_out417, gat_out424, gat_out425, gat_out426, gat_out427, gat_out432, gat_out437, gat_out442, gat_out443, gat_out444, gat_out445, gat_out451, gat_out460, gat_out463, gat_out466, gat_out475, gat_out476, gat_out477, gat_out478, gat_out479, gat_out480, gat_out481, gat_out482, gat_out483, gat_out488, gat_out489, gat_out490, gat_out491, gat_out492, gat_out495, gat_out498, gat_out499, gat_out500, gat_out501, gat_out502, gat_out503, gat_out504, gat_out505, gat_out506, gat_out507, gat_out508, gat_out509, gat_out510, gat_out511, gat_out512, gat_out513, gat_out514, gat_out515, gat_out516, gat_out517, gat_out518, gat_out519, gat_out520, gat_out521, gat_out522, gat_out523, gat_out524, gat_out525, gat_out526, gat_out527, gat_out528, gat_out529, gat_out530, gat_out533, gat_out536, gat_out537, gat_out538, gat_out539, gat_out540, gat_out541, gat_out542, gat_out543, gat_out544, gat_out547, gat_out550, gat_out551, gat_out552, gat_out553, gat_out557, gat_out561, gat_out565, gat_out569, gat_out573, gat_out577, gat_out581, gat_out585, gat_out586, gat_out587, gat_out588, gat_out589, gat_out590, gat_out593, gat_out596, gat_out597, gat_out600, gat_out605, gat_out606, gat_out609, gat_out615, gat_out616, gat_out619, gat_out624, gat_out625, gat_out628, gat_out631, gat_out632, gat_out635, gat_out640, gat_out641, gat_out644, gat_out650, gat_out651, gat_out654, gat_out659, gat_out660, gat_out661, gat_out662, gat_out665, gat_out669, gat_out670, gat_out673, gat_out677, gat_out678, gat_out682, gat_out686, gat_out687, gat_out692, gat_out696, gat_out697, gat_out700, gat_out704, gat_out705, gat_out708, gat_out712, gat_out713, gat_out717, gat_out721, gat_out722, gat_out727, gat_out731, gat_out732, gat_out733, gat_out734, gat_out735, gat_out736, gat_out737, gat_out738, gat_out739, gat_out740, gat_out741, gat_out742, gat_out743, gat_out744, gat_out745, gat_out746, gat_out747, gat_out748, gat_out749, gat_out750, gat_out751, gat_out752, gat_out753, gat_out754, gat_out755, gat_out756, gat_out757, gat_out758, gat_out759, gat_out760, gat_out761, gat_out762, gat_out763, gat_out764, gat_out765, gat_out766, gat_out769, gat_out770, gat_out771, gat_out772, gat_out773, gat_out777, gat_out778, gat_out781, gat_out782, gat_out785, gat_out786, gat_out787, gat_out788, gat_out789, gat_out790, gat_out791, gat_out792, gat_out793, gat_out794, gat_out795, gat_out796, gat_out802, gat_out803, gat_out804, gat_out805, gat_out806, gat_out807, gat_out808, gat_out809, gat_out810, gat_out811, gat_out812, gat_out813, gat_out814, gat_out815, gat_out819, gat_out822, gat_out825, gat_out826, gat_out827, gat_out828, gat_out829, gat_out830, gat_out831, gat_out832, gat_out833, gat_out834, gat_out835, gat_out836, gat_out837, gat_out838, gat_out839, gat_out840, gat_out841, gat_out842, gat_out843, gat_out844, gat_out845, gat_out846, gat_out847, gat_out848, gat_out849, gat_out851, gat_out852, gat_out853, gat_out854, gat_out855, gat_out856, gat_out857, gat_out858, gat_out859, gat_out860, gat_out861, gat_out862, gat_out867, gat_out868, gat_out869, gat_out870, gat_out871, gat_out872, gat_out873, gat_out875, gat_out876, gat_out877;
nand gat269 (gat_out269, gat1, gat8, gat13, gat17);
nand gat270 (gat_out270, gat1, gat26, gat13, gat17);
and gat273 (gat_out273, gat29, gat36, gat42);
and gat276 (gat_out276, gat1, gat26, gat51);
nand gat279 (gat_out279, gat1, gat8, gat51, gat17);
nand gat280 (gat_out280, gat1, gat8, gat13, gat55);
nand gat284 (gat_out284, gat59, gat42, gat68, gat72);
nand gat285 (gat_out285, gat29, gat68);
nand gat286 (gat_out286, gat59, gat68, gat74);
and gat287 (gat_out287, gat29, gat75, gat80);
and gat290 (gat_out290, gat29, gat75, gat42);
and gat291 (gat_out291, gat29, gat36, gat80);
and gat292 (gat_out292, gat29, gat36, gat42);
and gat293 (gat_out293, gat59, gat75, gat80);
and gat294 (gat_out294, gat59, gat75, gat42);
and gat295 (gat_out295, gat59, gat36, gat80);
and gat296 (gat_out296, gat59, gat36, gat42);
and gat297 (gat_out297, gat85, gat86);
or gat298 (gat_out298, gat87, gat88);
nand gat301 (gat_out301, gat91, gat96);
or gat302 (gat_out302, gat91, gat96);
nand gat303 (gat_out303, gat101, gat106);
or gat304 (gat_out304, gat101, gat106);
nand gat305 (gat_out305, gat111, gat116);
or gat306 (gat_out306, gat111, gat116);
nand gat307 (gat_out307, gat121, gat126);
or gat308 (gat_out308, gat121, gat126);
and gat309 (gat_out309, gat8, gat138);
not gat310 (gat_out310, gat268);
and gat316 (gat_out316, gat51, gat138);
and gat317 (gat_out317, gat17, gat138);
and gat318 (gat_out318, gat152, gat138);
nand gat319 (gat_out319, gat59, gat156);
nor gat322 (gat_out322, gat17, gat42);
and gat323 (gat_out323, gat17, gat42);
nand gat324 (gat_out324, gat159, gat165);
or gat325 (gat_out325, gat159, gat165);
nand gat326 (gat_out326, gat171, gat177);
or gat327 (gat_out327, gat171, gat177);
nand gat328 (gat_out328, gat183, gat189);
or gat329 (gat_out329, gat183, gat189);
nand gat330 (gat_out330, gat195, gat201);
or gat331 (gat_out331, gat195, gat201);
and gat332 (gat_out332, gat210, gat91);
and gat333 (gat_out333, gat210, gat96);
and gat334 (gat_out334, gat210, gat101);
and gat335 (gat_out335, gat210, gat106);
and gat336 (gat_out336, gat210, gat111);
and gat337 (gat_out337, gat255, gat259);
and gat338 (gat_out338, gat210, gat116);
and gat339 (gat_out339, gat255, gat260);
and gat340 (gat_out340, gat210, gat121);
and gat341 (gat_out341, gat255, gat267);
not gat342 (gat_out342, gat_out269);
not gat343 (gat_out343, gat_out273);
or gat344 (gat_out344, gat_out270, gat_out273);
not gat345 (gat_out345, gat_out276);
not gat346 (gat_out346, gat_out276);
not gat347 (gat_out347, gat_out279);
nor gat348 (gat_out348, gat_out280, gat_out284);
or gat349 (gat_out349, gat_out280, gat_out285);
or gat350 (gat_out350, gat_out280, gat_out286);
not gat351 (gat_out351, gat_out293);
not gat352 (gat_out352, gat_out294);
not gat353 (gat_out353, gat_out295);
not gat354 (gat_out354, gat_out296);
nand gat355 (gat_out355, gat89, gat_out298);
and gat356 (gat_out356, gat90, gat_out298);
nand gat357 (gat_out357, gat_out301, gat_out302);
nand gat360 (gat_out360, gat_out303, gat_out304);
nand gat363 (gat_out363, gat_out305, gat_out306);
nand gat366 (gat_out366, gat_out307, gat_out308);
not gat369 (gat_out369, gat_out310);
nor gat375 (gat_out375, gat_out322, gat_out323);
nand gat376 (gat_out376, gat_out324, gat_out325);
nand gat379 (gat_out379, gat_out326, gat_out327);
nand gat382 (gat_out382, gat_out328, gat_out329);
nand gat385 (gat_out385, gat_out330, gat_out331);
buf gat388 (gat_out388, gat_out290);
buf gat389 (gat_out389, gat_out291);
buf gat390 (gat_out390, gat_out292);
buf gat391 (gat_out391, gat_out297);
or gat392 (gat_out392, gat_out270, gat_out343);
not gat393 (gat_out393, gat_out345);
not gat399 (gat_out399, gat_out346);
and gat400 (gat_out400, gat_out348, gat73);
not gat401 (gat_out401, gat_out349);
not gat402 (gat_out402, gat_out350);
not gat403 (gat_out403, gat_out355);
not gat404 (gat_out404, gat_out357);
not gat405 (gat_out405, gat_out360);
and gat406 (gat_out406, gat_out357, gat_out360);
not gat407 (gat_out407, gat_out363);
not gat408 (gat_out408, gat_out366);
and gat409 (gat_out409, gat_out363, gat_out366);
nand gat410 (gat_out410, gat_out347, gat_out352);
not gat411 (gat_out411, gat_out376);
not gat412 (gat_out412, gat_out379);
and gat413 (gat_out413, gat_out376, gat_out379);
not gat414 (gat_out414, gat_out382);
not gat415 (gat_out415, gat_out385);
and gat416 (gat_out416, gat_out382, gat_out385);
and gat417 (gat_out417, gat210, gat_out369);
buf gat418 (gat_out418, gat_out342);
buf gat419 (gat_out419, gat_out344);
buf gat420 (gat_out420, gat_out351);
buf gat421 (gat_out421, gat_out353);
buf gat422 (gat_out422, gat_out354);
buf gat423 (gat_out423, gat_out356);
not gat424 (gat_out424, gat_out400);
and gat425 (gat_out425, gat_out404, gat_out405);
and gat426 (gat_out426, gat_out407, gat_out408);
and gat427 (gat_out427, gat_out319, gat_out393, gat55);
and gat432 (gat_out432, gat_out393, gat17, gat_out287);
nand gat437 (gat_out437, gat_out393, gat_out287, gat55);
nand gat442 (gat_out442, gat_out375, gat59, gat156, gat_out393);
nand gat443 (gat_out443, gat_out393, gat_out319, gat17);
and gat444 (gat_out444, gat_out411, gat_out412);
and gat445 (gat_out445, gat_out414, gat_out415);
buf gat446 (gat_out446, gat_out392);
buf gat447 (gat_out447, gat_out399);
buf gat448 (gat_out448, gat_out401);
buf gat449 (gat_out449, gat_out402);
buf gat450 (gat_out450, gat_out403);
not gat451 (gat_out451, gat_out424);
nor gat460 (gat_out460, gat_out406, gat_out425);
nor gat463 (gat_out463, gat_out409, gat_out426);
nand gat466 (gat_out466, gat_out442, gat_out410);
and gat475 (gat_out475, gat143, gat_out427);
and gat476 (gat_out476, gat_out310, gat_out432);
and gat477 (gat_out477, gat146, gat_out427);
and gat478 (gat_out478, gat_out310, gat_out432);
and gat479 (gat_out479, gat149, gat_out427);
and gat480 (gat_out480, gat_out310, gat_out432);
and gat481 (gat_out481, gat153, gat_out427);
and gat482 (gat_out482, gat_out310, gat_out432);
nand gat483 (gat_out483, gat_out443, gat1);
or gat488 (gat_out488, gat_out369, gat_out437);
or gat489 (gat_out489, gat_out369, gat_out437);
or gat490 (gat_out490, gat_out369, gat_out437);
or gat491 (gat_out491, gat_out369, gat_out437);
nor gat492 (gat_out492, gat_out413, gat_out444);
nor gat495 (gat_out495, gat_out416, gat_out445);
nand gat498 (gat_out498, gat130, gat_out460);
or gat499 (gat_out499, gat130, gat_out460);
nand gat500 (gat_out500, gat_out463, gat135);
or gat501 (gat_out501, gat_out463, gat135);
and gat502 (gat_out502, gat91, gat_out466);
nor gat503 (gat_out503, gat_out475, gat_out476);
and gat504 (gat_out504, gat96, gat_out466);
nor gat505 (gat_out505, gat_out477, gat_out478);
and gat506 (gat_out506, gat101, gat_out466);
nor gat507 (gat_out507, gat_out479, gat_out480);
and gat508 (gat_out508, gat106, gat_out466);
nor gat509 (gat_out509, gat_out481, gat_out482);
and gat510 (gat_out510, gat143, gat_out483);
and gat511 (gat_out511, gat111, gat_out466);
and gat512 (gat_out512, gat146, gat_out483);
and gat513 (gat_out513, gat116, gat_out466);
and gat514 (gat_out514, gat149, gat_out483);
and gat515 (gat_out515, gat121, gat_out466);
and gat516 (gat_out516, gat153, gat_out483);
and gat517 (gat_out517, gat126, gat_out466);
nand gat518 (gat_out518, gat130, gat_out492);
or gat519 (gat_out519, gat130, gat_out492);
nand gat520 (gat_out520, gat_out495, gat207);
or gat521 (gat_out521, gat_out495, gat207);
and gat522 (gat_out522, gat_out451, gat159);
and gat523 (gat_out523, gat_out451, gat165);
and gat524 (gat_out524, gat_out451, gat171);
and gat525 (gat_out525, gat_out451, gat177);
and gat526 (gat_out526, gat_out451, gat183);
nand gat527 (gat_out527, gat_out451, gat189);
nand gat528 (gat_out528, gat_out451, gat195);
nand gat529 (gat_out529, gat_out451, gat201);
nand gat530 (gat_out530, gat_out498, gat_out499);
nand gat533 (gat_out533, gat_out500, gat_out501);
nor gat536 (gat_out536, gat_out309, gat_out502);
nor gat537 (gat_out537, gat_out316, gat_out504);
nor gat538 (gat_out538, gat_out317, gat_out506);
nor gat539 (gat_out539, gat_out318, gat_out508);
nor gat540 (gat_out540, gat_out510, gat_out511);
nor gat541 (gat_out541, gat_out512, gat_out513);
nor gat542 (gat_out542, gat_out514, gat_out515);
nor gat543 (gat_out543, gat_out516, gat_out517);
nand gat544 (gat_out544, gat_out518, gat_out519);
nand gat547 (gat_out547, gat_out520, gat_out521);
not gat550 (gat_out550, gat_out530);
not gat551 (gat_out551, gat_out533);
and gat552 (gat_out552, gat_out530, gat_out533);
nand gat553 (gat_out553, gat_out536, gat_out503);
nand gat557 (gat_out557, gat_out537, gat_out505);
nand gat561 (gat_out561, gat_out538, gat_out507);
nand gat565 (gat_out565, gat_out539, gat_out509);
nand gat569 (gat_out569, gat_out488, gat_out540);
nand gat573 (gat_out573, gat_out489, gat_out541);
nand gat577 (gat_out577, gat_out490, gat_out542);
nand gat581 (gat_out581, gat_out491, gat_out543);
not gat585 (gat_out585, gat_out544);
not gat586 (gat_out586, gat_out547);
and gat587 (gat_out587, gat_out544, gat_out547);
and gat588 (gat_out588, gat_out550, gat_out551);
and gat589 (gat_out589, gat_out585, gat_out586);
nand gat590 (gat_out590, gat_out553, gat159);
or gat593 (gat_out593, gat_out553, gat159);
and gat596 (gat_out596, gat246, gat_out553);
nand gat597 (gat_out597, gat_out557, gat165);
or gat600 (gat_out600, gat_out557, gat165);
and gat605 (gat_out605, gat246, gat_out557);
nand gat606 (gat_out606, gat_out561, gat171);
or gat609 (gat_out609, gat_out561, gat171);
and gat615 (gat_out615, gat246, gat_out561);
nand gat616 (gat_out616, gat_out565, gat177);
or gat619 (gat_out619, gat_out565, gat177);
and gat624 (gat_out624, gat246, gat_out565);
nand gat625 (gat_out625, gat_out569, gat183);
or gat628 (gat_out628, gat_out569, gat183);
and gat631 (gat_out631, gat246, gat_out569);
nand gat632 (gat_out632, gat_out573, gat189);
or gat635 (gat_out635, gat_out573, gat189);
and gat640 (gat_out640, gat246, gat_out573);
nand gat641 (gat_out641, gat_out577, gat195);
or gat644 (gat_out644, gat_out577, gat195);
and gat650 (gat_out650, gat246, gat_out577);
nand gat651 (gat_out651, gat_out581, gat201);
or gat654 (gat_out654, gat_out581, gat201);
and gat659 (gat_out659, gat246, gat_out581);
nor gat660 (gat_out660, gat_out552, gat_out588);
nor gat661 (gat_out661, gat_out587, gat_out589);
not gat662 (gat_out662, gat_out590);
and gat665 (gat_out665, gat_out593, gat_out590);
nor gat669 (gat_out669, gat_out596, gat_out522);
not gat670 (gat_out670, gat_out597);
and gat673 (gat_out673, gat_out600, gat_out597);
nor gat677 (gat_out677, gat_out605, gat_out523);
not gat678 (gat_out678, gat_out606);
and gat682 (gat_out682, gat_out609, gat_out606);
nor gat686 (gat_out686, gat_out615, gat_out524);
not gat687 (gat_out687, gat_out616);
and gat692 (gat_out692, gat_out619, gat_out616);
nor gat696 (gat_out696, gat_out624, gat_out525);
not gat697 (gat_out697, gat_out625);
and gat700 (gat_out700, gat_out628, gat_out625);
nor gat704 (gat_out704, gat_out631, gat_out526);
not gat705 (gat_out705, gat_out632);
and gat708 (gat_out708, gat_out635, gat_out632);
nor gat712 (gat_out712, gat_out337, gat_out640);
not gat713 (gat_out713, gat_out641);
and gat717 (gat_out717, gat_out644, gat_out641);
nor gat721 (gat_out721, gat_out339, gat_out650);
not gat722 (gat_out722, gat_out651);
and gat727 (gat_out727, gat_out654, gat_out651);
nor gat731 (gat_out731, gat_out341, gat_out659);
nand gat732 (gat_out732, gat_out654, gat261);
nand gat733 (gat_out733, gat_out644, gat_out654, gat261);
nand gat734 (gat_out734, gat_out635, gat_out644, gat_out654, gat261);
not gat735 (gat_out735, gat_out662);
and gat736 (gat_out736, gat228, gat_out665);
and gat737 (gat_out737, gat237, gat_out662);
not gat738 (gat_out738, gat_out670);
and gat739 (gat_out739, gat228, gat_out673);
and gat740 (gat_out740, gat237, gat_out670);
not gat741 (gat_out741, gat_out678);
and gat742 (gat_out742, gat228, gat_out682);
and gat743 (gat_out743, gat237, gat_out678);
not gat744 (gat_out744, gat_out687);
and gat745 (gat_out745, gat228, gat_out692);
and gat746 (gat_out746, gat237, gat_out687);
not gat747 (gat_out747, gat_out697);
and gat748 (gat_out748, gat228, gat_out700);
and gat749 (gat_out749, gat237, gat_out697);
not gat750 (gat_out750, gat_out705);
and gat751 (gat_out751, gat228, gat_out708);
and gat752 (gat_out752, gat237, gat_out705);
not gat753 (gat_out753, gat_out713);
and gat754 (gat_out754, gat228, gat_out717);
and gat755 (gat_out755, gat237, gat_out713);
not gat756 (gat_out756, gat_out722);
nor gat757 (gat_out757, gat_out727, gat261);
and gat758 (gat_out758, gat_out727, gat261);
and gat759 (gat_out759, gat228, gat_out727);
and gat760 (gat_out760, gat237, gat_out722);
nand gat761 (gat_out761, gat_out644, gat_out722);
nand gat762 (gat_out762, gat_out635, gat_out713);
nand gat763 (gat_out763, gat_out635, gat_out644, gat_out722);
nand gat764 (gat_out764, gat_out609, gat_out687);
nand gat765 (gat_out765, gat_out600, gat_out678);
nand gat766 (gat_out766, gat_out600, gat_out609, gat_out687);
buf gat767 (gat_out767, gat_out660);
buf gat768 (gat_out768, gat_out661);
nor gat769 (gat_out769, gat_out736, gat_out737);
nor gat770 (gat_out770, gat_out739, gat_out740);
nor gat771 (gat_out771, gat_out742, gat_out743);
nor gat772 (gat_out772, gat_out745, gat_out746);
nand gat773 (gat_out773, gat_out750, gat_out762, gat_out763, gat_out734);
nor gat777 (gat_out777, gat_out748, gat_out749);
nand gat778 (gat_out778, gat_out753, gat_out761, gat_out733);
nor gat781 (gat_out781, gat_out751, gat_out752);
nand gat782 (gat_out782, gat_out756, gat_out732);
nor gat785 (gat_out785, gat_out754, gat_out755);
nor gat786 (gat_out786, gat_out757, gat_out758);
nor gat787 (gat_out787, gat_out759, gat_out760);
nor gat788 (gat_out788, gat_out700, gat_out773);
and gat789 (gat_out789, gat_out700, gat_out773);
nor gat790 (gat_out790, gat_out708, gat_out778);
and gat791 (gat_out791, gat_out708, gat_out778);
nor gat792 (gat_out792, gat_out717, gat_out782);
and gat793 (gat_out793, gat_out717, gat_out782);
and gat794 (gat_out794, gat219, gat_out786);
nand gat795 (gat_out795, gat_out628, gat_out773);
nand gat796 (gat_out796, gat_out795, gat_out747);
nor gat802 (gat_out802, gat_out788, gat_out789);
nor gat803 (gat_out803, gat_out790, gat_out791);
nor gat804 (gat_out804, gat_out792, gat_out793);
nor gat805 (gat_out805, gat_out340, gat_out794);
nor gat806 (gat_out806, gat_out692, gat_out796);
and gat807 (gat_out807, gat_out692, gat_out796);
and gat808 (gat_out808, gat219, gat_out802);
and gat809 (gat_out809, gat219, gat_out803);
and gat810 (gat_out810, gat219, gat_out804);
nand gat811 (gat_out811, gat_out805, gat_out787, gat_out731, gat_out529);
nand gat812 (gat_out812, gat_out619, gat_out796);
nand gat813 (gat_out813, gat_out609, gat_out619, gat_out796);
nand gat814 (gat_out814, gat_out600, gat_out609, gat_out619, gat_out796);
nand gat815 (gat_out815, gat_out738, gat_out765, gat_out766, gat_out814);
nand gat819 (gat_out819, gat_out741, gat_out764, gat_out813);
nand gat822 (gat_out822, gat_out744, gat_out812);
nor gat825 (gat_out825, gat_out806, gat_out807);
nor gat826 (gat_out826, gat_out335, gat_out808);
nor gat827 (gat_out827, gat_out336, gat_out809);
nor gat828 (gat_out828, gat_out338, gat_out810);
not gat829 (gat_out829, gat_out811);
nor gat830 (gat_out830, gat_out665, gat_out815);
and gat831 (gat_out831, gat_out665, gat_out815);
nor gat832 (gat_out832, gat_out673, gat_out819);
and gat833 (gat_out833, gat_out673, gat_out819);
nor gat834 (gat_out834, gat_out682, gat_out822);
and gat835 (gat_out835, gat_out682, gat_out822);
and gat836 (gat_out836, gat219, gat_out825);
nand gat837 (gat_out837, gat_out826, gat_out777, gat_out704);
nand gat838 (gat_out838, gat_out827, gat_out781, gat_out712, gat_out527);
nand gat839 (gat_out839, gat_out828, gat_out785, gat_out721, gat_out528);
not gat840 (gat_out840, gat_out829);
nand gat841 (gat_out841, gat_out815, gat_out593);
nor gat842 (gat_out842, gat_out830, gat_out831);
nor gat843 (gat_out843, gat_out832, gat_out833);
nor gat844 (gat_out844, gat_out834, gat_out835);
nor gat845 (gat_out845, gat_out334, gat_out836);
not gat846 (gat_out846, gat_out837);
not gat847 (gat_out847, gat_out838);
not gat848 (gat_out848, gat_out839);
and gat849 (gat_out849, gat_out735, gat_out841);
buf gat850 (gat_out850, gat_out840);
and gat851 (gat_out851, gat219, gat_out842);
and gat852 (gat_out852, gat219, gat_out843);
and gat853 (gat_out853, gat219, gat_out844);
nand gat854 (gat_out854, gat_out845, gat_out772, gat_out696);
not gat855 (gat_out855, gat_out846);
not gat856 (gat_out856, gat_out847);
not gat857 (gat_out857, gat_out848);
not gat858 (gat_out858, gat_out849);
nor gat859 (gat_out859, gat_out417, gat_out851);
nor gat860 (gat_out860, gat_out332, gat_out852);
nor gat861 (gat_out861, gat_out333, gat_out853);
not gat862 (gat_out862, gat_out854);
buf gat863 (gat_out863, gat_out855);
buf gat864 (gat_out864, gat_out856);
buf gat865 (gat_out865, gat_out857);
buf gat866 (gat_out866, gat_out858);
nand gat867 (gat_out867, gat_out859, gat_out769, gat_out669);
nand gat868 (gat_out868, gat_out860, gat_out770, gat_out677);
nand gat869 (gat_out869, gat_out861, gat_out771, gat_out686);
not gat870 (gat_out870, gat_out862);
not gat871 (gat_out871, gat_out867);
not gat872 (gat_out872, gat_out868);
not gat873 (gat_out873, gat_out869);
buf gat874 (gat_out874, gat_out870);
not gat875 (gat_out875, gat_out871);
not gat876 (gat_out876, gat_out872);
not gat877 (gat_out877, gat_out873);
buf gat878 (gat_out878, gat_out875);
buf gat879 (gat_out879, gat_out876);
buf gat880 (gat_out880, gat_out877);
endmodule